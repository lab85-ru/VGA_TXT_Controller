//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW1NZ-LV1FN32C6/I5
//Device: GW1NZ-1
//Created Time: Fri May 26 19:05:23 2023

module rom (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b1;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h000008CEEEEC0000000EFF73FFBFE000000E119D1151E0000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000008CC80000000000C88EFFEC80000000C88777CC80000000008CEC800000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0008CCCC82AEE000FFFFF39DD93FFFFF00000C6226C00000FFFFFF7337FFFFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'h000088BC7CB880000006773333F3F0000000000000F3F00000088E8C6666C000;
defparam prom_inst_0.INIT_RAM_04 = 256'h000660666666600000008CE888EC800000026EEEEEEE620000000008E8000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h000E8CE888EC8000000EEEE000000000000C6C8C66C806C0000BBBBBBBBBF000;
defparam prom_inst_0.INIT_RAM_06 = 256'h00000000E00000000000008CEC8000000008CE88888880000008888888EC8000;
defparam prom_inst_0.INIT_RAM_07 = 256'h00000088CCEE000000000EECC88000000000008CEC800000000000E000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h000CCECCCECC00000000000000046660000880888CCC80000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h00000000000000000006CCCC68CC800000066008C6200000088C6666C026C880;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000088E88000000000006CFC600000000008CCCCCC80000000C80000008C000;
defparam prom_inst_0.INIT_RAM_0B = 256'h00000008C620000000088000000000000000000E000000000088800000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h000C6666C666C000000E60008C66C000000E8888888880000008C666666C8000;
defparam prom_inst_0.INIT_RAM_0D = 256'h00000008C666E000000C6666C0008000000C6666C000E000000ECCCECCCCC000;
defparam prom_inst_0.INIT_RAM_0E = 256'h000880008800000000088000880000000008C666E666C000000C6666C666C000;
defparam prom_inst_0.INIT_RAM_0F = 256'h000880888C66C000000008C6C8000000000000E00E0000000006C80008C60000;
defparam prom_inst_0.INIT_RAM_10 = 256'h000C62000026C000000C6666C666C0000006666E66C80000000C0CEEE66C0000;
defparam prom_inst_0.INIT_RAM_11 = 256'h000A666E0026C000000000088826E000000E62088826E0000008C666666C8000;
defparam prom_inst_0.INIT_RAM_12 = 256'h000666C88C6660000008CCCCCCCCE000000C88888888C00000066666E6666000;
defparam prom_inst_0.INIT_RAM_13 = 256'h000C66666666C0000006666EEE666000000666666EEE6000000E620000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h000C666C8066C0000006666CC666C0000ECCE6666666C00000000000C666C000;
defparam prom_inst_0.INIT_RAM_15 = 256'h000CEE666666600000008C6666666000000C666666666000000C888888AEE000;
defparam prom_inst_0.INIT_RAM_16 = 256'h000C00000000C000000E62008C66E000000C8888C666600000066CC88CC66000;
defparam prom_inst_0.INIT_RAM_17 = 256'h00F000000000000000000000000000C8000CCCCCCCCCC00000026EC800000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h000C60006C000000000C6666C80000000006CCCCC80000000000000000000080;
defparam prom_inst_0.INIT_RAM_19 = 256'h8CCCCCCCC6000000000800008026C000000C600E6C0000000006CCCCCCCCC000;
defparam prom_inst_0.INIT_RAM_1A = 256'h00066C88C6000000C66666666E066000000C888888088000000666666C000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h000C66666C000000000666666C00000000066666EC000000000C888888888000;
defparam prom_inst_0.INIT_RAM_1C = 256'h000C6C806C000000000000066C000000ECCCCCCCC6000000000C66666C000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h000CE666660000000008C666660000000006CCCCCC000000000C60000C000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h000E88880888E000000E6008CE0000008C6E6666660000000006C888C6000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h000E666C8000000000000000000000C600008888E88800000008888888888000;
defparam prom_inst_0.INIT_RAM_20 = 256'h000000002E08C6000888000000000000000000000026E08C000C6666C000C000;
defparam prom_inst_0.INIT_RAM_21 = 256'h00088EE88EE88000000888888EE88000000BB0000000000084CC000000000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h0008000800000000000CAAAAC888C000000BB0008C620000000C60000806C000;
defparam prom_inst_0.INIT_RAM_23 = 256'h000ECCCCCCCCE00000066666C000C00000066CC88CC6608C000CAAAAC8888000;
defparam prom_inst_0.INIT_RAM_24 = 256'h000000000000CC84000000000000088800000000000088080C66666C00800000;
defparam prom_inst_0.INIT_RAM_25 = 256'h0000000F000000000000000E000000000000000CEEEC000000000000000084CC;
defparam prom_inst_0.INIT_RAM_26 = 256'h00008C8000000000000CAAAC8C0000000000000005FB10000000000000000000;
defparam prom_inst_0.INIT_RAM_27 = 256'h000ECCCCCE00000000066666C008000000066C88C608C600000CAAAC88000000;
defparam prom_inst_0.INIT_RAM_28 = 256'h0008CCCCCCCCE000C66E6666660C6000000C666E666660C60000000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h000C6C8C66C806C00008888800888880000000000000E6200006C6666C600000;
defparam prom_inst_0.INIT_RAM_2A = 256'h0006C8C600000000000C60088806C000000C2A2222A2C000000E62088826E0C0;
defparam prom_inst_0.INIT_RAM_2B = 256'h000C88888888C060000C2AA2AA22C0000000000E00000000000006666E000000;
defparam prom_inst_0.INIT_RAM_2C = 256'h000C888888080000000C88888888C0000000E0088E8800000000000008CC8000;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000000800000000000BBBBBBBBBF000000C666666000000000000000E220000;
defparam prom_inst_0.INIT_RAM_2E = 256'h0008C6C800000000000C60806C000000000CCCCCFCFDF000000C60C66C0C0000;
defparam prom_inst_0.INIT_RAM_2F = 256'h000C8888880C0000000C6C806C000000000C666C8066C000C66666666E066000;
defparam prom_inst_0.INIT_RAM_30 = 256'h000000000026E000000C6666C666C000000C6666C002E0000006666E6666E000;
defparam prom_inst_0.INIT_RAM_31 = 256'h000C6666C666C0000006644CC4466000000E62088826E000013F66666666E000;
defparam prom_inst_0.INIT_RAM_32 = 256'h000666666666E00000066CC88CC6600000066666EE6660C600066666EE666000;
defparam prom_inst_0.INIT_RAM_33 = 256'h000666666666E000000C66666666C00000066666E6666000000666666EEE6000;
defparam prom_inst_0.INIT_RAM_34 = 256'h000C666E66666000000C888888AEE000000C62000066C0000000000C6666C000;
defparam prom_inst_0.INIT_RAM_35 = 256'h0006666E66666000033F66666666600000066CC88CC6600000080C666666C000;
defparam prom_inst_0.INIT_RAM_36 = 256'h0006EEEE66666000000C6666C0008000033F666666666000000E666666666000;
defparam prom_inst_0.INIT_RAM_37 = 256'h000ECCCCCCCCE000000C66666666C000000C6666E666C000000C6666C0000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h000000022E000000000C66C66C000000000C6666C00C60000006CCCCC8000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h000C66C66C000000000664C466000000000C60E66C000000033F66666E000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h000666666E00000000066C88C6000000000666EE660C6000000666EE66000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h000666666E000000000C66666C000000000666E666000000000666EEE6000000;
defparam prom_inst_0.INIT_RAM_3C = 256'hC66E666666000000000C8888AE000000000C60006C000000000C66666C000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h00066E6666000000033F6666660000000006C888C6000000800C66666C080000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0006EE6666000000000C66C008000000033E666666000000000E666666000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h000ECCCCCE000000000C66666C000000000C66E66C000000000C66C000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b1;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0000137FFFF600000007FFECFFDF70000007889B88A870000000000000000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h000000133100000000003117FF7310000000311EEE33100000000137F7310000;
defparam prom_inst_1.INIT_RAM_02 = 256'h0007CCCC73101000FFFFFC9BB9CFFFFF0000036446300000FFFFFFECCEFFFFFF;
defparam prom_inst_1.INIT_RAM_03 = 256'h000011D3E3D1100000CEE66666767000000EF733333330000001171366663000;
defparam prom_inst_1.INIT_RAM_04 = 256'h0006606666666000000013711173100000000013F31000000008CEFFFFFEC800;
defparam prom_inst_1.INIT_RAM_05 = 256'h0007137111731000000FFFF0000000000007C036CC636C70000111117DDD7000;
defparam prom_inst_1.INIT_RAM_06 = 256'h00000036F630000000000010F010000000013711111110000001111111731000;
defparam prom_inst_1.INIT_RAM_07 = 256'h0000013377FF000000000FF77331000000000026F6200000000000FCCC000000;
defparam prom_inst_1.INIT_RAM_08 = 256'h00066F666F660000000000000002666000011011133310000000000000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h00000000063330000007CCCD736630000008C6310CC000000117C8007CCC7110;
defparam prom_inst_1.INIT_RAM_0A = 256'h00000117110000000000063F3600000000031000000130000000133333310000;
defparam prom_inst_1.INIT_RAM_0B = 256'h0008C6310000000000011000000000000000000F000000000311100000000000;
defparam prom_inst_1.INIT_RAM_0C = 256'h0007C000300C7000000FCC63100C7000000711111173100000036CCDDCC63000;
defparam prom_inst_1.INIT_RAM_0D = 256'h00033331000CF0000007CCCCFCC630000007C000FCCCF0000001000FC6310000;
defparam prom_inst_1.INIT_RAM_0E = 256'h00311000110000000001100011000000000700007CCC70000007CCCC7CCC7000;
defparam prom_inst_1.INIT_RAM_0F = 256'h0001101110CC7000000631000136000000000070070000000000013631000000;
defparam prom_inst_1.INIT_RAM_10 = 256'h00036CCCCCC63000000F66667666F000000CCCCFCC6310000007CDDDDCC70000;
defparam prom_inst_1.INIT_RAM_11 = 256'h00036CCDCCC63000000F66667666F000000F66667666F000000F66666666F000;
defparam prom_inst_1.INIT_RAM_12 = 256'h000E66677666E0000007CCC0000010000003111111113000000CCCCCFCCCC000;
defparam prom_inst_1.INIT_RAM_13 = 256'h0007CCCCCCCC7000000CCCCCDFFEC000000CCCCCDFFEC000000F66666666F000;
defparam prom_inst_1.INIT_RAM_14 = 256'h0007CC0036CC7000000E66667666F0000007DDCCCCCC7000000F66667666F000;
defparam prom_inst_1.INIT_RAM_15 = 256'h0006EFDDDCCCC000000136CCCCCCC0000007CCCCCCCCC0000003111111577000;
defparam prom_inst_1.INIT_RAM_16 = 256'h0003333333333000000FCC63108CF0000003111136666000000CC673376CC000;
defparam prom_inst_1.INIT_RAM_17 = 256'h00F000000000000000000000000000630003000000003000000000137EC80000;
defparam prom_inst_1.INIT_RAM_18 = 256'h0007CCCCC7000000000766666766E0000007CCC7070000000000000000000013;
defparam prom_inst_1.INIT_RAM_19 = 256'h7C07CCCCC700000000073333733310000007CCCFC70000000007CCCC63001000;
defparam prom_inst_1.INIT_RAM_1A = 256'h000E66776666E00036600000000000000003111113011000000E66667666E000;
defparam prom_inst_1.INIT_RAM_1B = 256'h0007CCCCC7000000000666666D000000000CDDDDFE0000000003111111113000;
defparam prom_inst_1.INIT_RAM_1C = 256'h0007C036C7000000000F66667D0000001007CCCCC7000000F66766666D000000;
defparam prom_inst_1.INIT_RAM_1D = 256'h0006FDDDCC00000000036CCCCC0000000007CCCCCC000000000133333F331000;
defparam prom_inst_1.INIT_RAM_1E = 256'h0000111171110000000FC631CF000000F007CCCCCC000000000C63336C000000;
defparam prom_inst_1.INIT_RAM_1F = 256'h000FCCC63100000000000000000000D700071111011170000001111111111000;
defparam prom_inst_1.INIT_RAM_20 = 256'h000F66666F0100001011000000000000000F66666666F010000E66676666F000;
defparam prom_inst_1.INIT_RAM_21 = 256'h00011771177110000001111117711000000DD000000000004266000000000000;
defparam prom_inst_1.INIT_RAM_22 = 256'h0001363100000000000D55555555F00000019C6310CC000000036CCFCFC63000;
defparam prom_inst_1.INIT_RAM_23 = 256'h001F66666666E000000E66667666F000000E66677666E010000DDDDDFDDDD000;
defparam prom_inst_1.INIT_RAM_24 = 256'h000000000000664200000000000010110000000000001110010E666766F66000;
defparam prom_inst_1.INIT_RAM_25 = 256'h0000000F000000000000000F0000000000000003777300000000000000004266;
defparam prom_inst_1.INIT_RAM_26 = 256'h0003101300000000000D55555F000000000000000555F0000000000000000000;
defparam prom_inst_1.INIT_RAM_27 = 256'h001F66666E000000000E6666766F6000000E66776E010000000DDDDFDD000000;
defparam prom_inst_1.INIT_RAM_28 = 256'h0007CCC0000010007C07CCCCCC07C0000007C007CCCCC07C0000000000000000;
defparam prom_inst_1.INIT_RAM_29 = 256'h0007C036CC636C700001111100111110000F66666666F000000C7CCCC7C00000;
defparam prom_inst_1.INIT_RAM_2A = 256'h00036D63000000000007CCCCFCCC7000000789AAAA987000000F66667666F060;
defparam prom_inst_1.INIT_RAM_2B = 256'h000311111111306000078AABAAB870000000000F00000000000000000F000000;
defparam prom_inst_1.INIT_RAM_2C = 256'h0003111113010000000311111111300000007001171100000000000003663000;
defparam prom_inst_1.INIT_RAM_2D = 256'h0000000100000000000111117DDD7000C667666666000000000F66666F000000;
defparam prom_inst_1.INIT_RAM_2E = 256'h000D636D000000000007CCFCC7000000000CCCDDFEECC0000007CCFCC7060000;
defparam prom_inst_1.INIT_RAM_2F = 256'h00031111130600000007C036C70000000007CC0036CC70003660000000000000;
defparam prom_inst_1.INIT_RAM_30 = 256'h000F66666666F000000F66667666F000000F66667666F000000CCCCFCC631000;
defparam prom_inst_1.INIT_RAM_31 = 256'h0007C000300C7000000DD557755DD000000F66667666F00008CF666666631000;
defparam prom_inst_1.INIT_RAM_32 = 256'h000C666666631000000E66677666E000000CCCEFDCCCC07C000CCCEFDCCCC000;
defparam prom_inst_1.INIT_RAM_33 = 256'h000CCCCCCCCCF0000007CCCCCCCC7000000CCCCCFCCCC000000CCCCCDFFEC000;
defparam prom_inst_1.INIT_RAM_34 = 256'h0007C007CCCCC00000031111115770000007CCCCCCCC7000000F66676666F000;
defparam prom_inst_1.INIT_RAM_35 = 256'h00000007CCCCC000000FCCCCCCCCC000000CC673376CC000000317DDDDDD7000;
defparam prom_inst_1.INIT_RAM_36 = 256'h000FDDDDFCCCC0000007333333BBF000000FDDDDDDDDD000000FDDDDDDDDD000;
defparam prom_inst_1.INIT_RAM_37 = 256'h000CCCC67CCC7000000CDDDDFDDDC0000007C002320C7000000F66667666F000;
defparam prom_inst_1.INIT_RAM_38 = 256'h000F66666F000000000F66766F0000000007CCCCFCC700000007CCC707000000;
defparam prom_inst_1.INIT_RAM_39 = 256'h0007C030C7000000000DD575DD0000000007CCFCC70000000CCF666631000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h000E666631000000000E66776E000000000CEFDCCC07C000000CEFDCCC000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h000CCCCCCF0000000007CCCCC7000000000CCCFCCC000000000CDDFFEC000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h7C07CCCCCC00000000031111570000000007CCCCC7000000F66766666D000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h000007CCCC000000000FCCCCCC000000000C63336C0000003117DDDDD7130000;
defparam prom_inst_1.INIT_RAM_3E = 256'h000FDDFCCC0000000007333BBF000000000FDDDDDD000000000FDDDDDD000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h000CC67CC7000000000CDDFDDC0000000007C030C7000000000F66766F000000;

endmodule //rom
