//`define VGA80x25 // font 8x16
//`define VGA64x30 // font 8x16

// set resolution
`define VGA80x25
//`define VGA64x30

// port intenal FPGA or SPI controller
//`define VGA_CMD_PORT

// port DMA for internal FPGA
//
`define VGA_DMA_PORT

